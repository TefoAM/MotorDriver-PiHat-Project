*SRC=1N4728A;DI_1N4728A;Diodes;Zener <=10V; 3.30V  1.00W   Diodes Inc.
Zener
*SYM=HZEN
.SUBCKT DI_1N4728A  1 2
*        Terminals    A   K
D1 1 2 DF
DZ 3 1 DR
VZ 2 3 0.972
.MODEL DF D ( IS=125p RS=0.620 N=1.10
+ CJO=364p VJ=0.750 M=0.330 TT=50.1n )
.MODEL DR D ( IS=25.0f RS=1.24 N=3.00 )
.ENDS